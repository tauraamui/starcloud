module data

fn test_matrix_init() {
	mat := Matrix.new(10, 5)
}
